//"interface.sv"

//Declare all the signals in interface use logic as datatype
interface intf();
  
  logic a;
  logic b;
  logic cin;
  logic s;
  logic cout;
  
endinterface

//No clocking and modport is not present here as this is not that complex design..
